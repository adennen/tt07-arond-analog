magic
tech sky130A
timestamp 1717269366
<< metal1 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -1100 5300 -100 6300 se
rect -100 5300 900 6300
tri -1600 4800 -1100 5300 se
tri -1100 4800 -600 5300 nw
tri -2100 4300 -1600 4800 se
tri -1600 4300 -1100 4800 nw
tri -2100 4157 -1957 4300 ne
rect -1957 4157 -1600 4300
tri -4207 3450 -3500 4157 se
tri -3500 3450 -2793 4157 sw
tri -1957 3800 -1600 4157 ne
tri -1600 3800 -1100 4300 sw
tri -4207 2743 -3500 3450 ne
tri -3500 2743 -2793 3450 nw
tri -1600 3300 -1100 3800 ne
tri -1100 3300 -600 3800 sw
rect -100 3300 400 5300
tri -1100 2743 -543 3300 ne
rect -543 2743 900 3300
tri -543 2300 -100 2743 ne
rect -100 2300 900 2743
rect -300 500 -100 700
tri -200 300 -100 400 se
tri -100 300 0 400 sw
rect 500 300 800 400
tri 800 300 900 400 sw
tri -300 200 -200 300 se
tri -200 200 -100 300 nw
tri -100 200 0 300 ne
tri 0 200 100 300 sw
tri -500 0 -300 200 se
tri -300 100 -200 200 nw
tri 0 100 100 200 ne
tri 100 100 200 200 sw
rect 100 0 200 100
tri 200 0 300 100 sw
rect -500 -100 300 0
rect -500 -200 -300 -100
rect 100 -200 300 -100
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal2 >>
rect -6100 18900 -5400 18950
rect -6300 18850 -5150 18900
rect -6500 18800 -5000 18850
rect -6600 18750 -4900 18800
rect -6700 18700 -4800 18750
rect -6800 18650 -4700 18700
rect -6900 18600 -4600 18650
rect -6950 18550 -4500 18600
rect -7050 18500 -4450 18550
rect -7100 18450 -4400 18500
rect -7150 18400 -4300 18450
rect -7250 18350 -4250 18400
rect -7300 18300 -4200 18350
rect -5450 18250 -4150 18300
rect -5500 18200 -4100 18250
rect -5500 18150 -4600 18200
rect -5550 18050 -4650 18150
rect -4550 18100 -4050 18200
rect -4550 18050 -4000 18100
rect -5600 17950 -4700 18050
rect -4550 18000 -3950 18050
rect -4550 17950 -3900 18000
rect -5650 17850 -4750 17950
rect -4500 17900 -3900 17950
rect -4500 17850 -3850 17900
rect -7700 17750 -6250 17800
rect -5700 17750 -4800 17850
rect -4500 17750 -3800 17850
rect -7750 17650 -6250 17750
rect -5750 17650 -4850 17750
rect -4500 17700 -3750 17750
rect -4450 17650 -3750 17700
rect -7800 17550 -6300 17650
rect -5800 17550 -4900 17650
rect -7850 17450 -6350 17550
rect -5850 17500 -4900 17550
rect -4450 17550 -3700 17650
rect -5850 17450 -4950 17500
rect -4450 17450 -3650 17550
rect -7850 17400 -6400 17450
rect -7900 17350 -6400 17400
rect -5900 17400 -4950 17450
rect -7900 17250 -6450 17350
rect -5900 17300 -5000 17400
rect -4400 17300 -3600 17450
rect -7950 17150 -6500 17250
rect -5950 17200 -5050 17300
rect -4400 17200 -3550 17300
rect -7950 17050 -6550 17150
rect -6000 17100 -5100 17200
rect -4350 17100 -3550 17200
rect -8000 16950 -6600 17050
rect -6050 17000 -5150 17100
rect -8000 16800 -6650 16950
rect -6100 16900 -5200 17000
rect -4350 16950 -3500 17100
rect -6150 16800 -5250 16900
rect -8000 16700 -6700 16800
rect -6200 16700 -5300 16800
rect -4800 16750 -4700 16850
rect -8000 16600 -6750 16700
rect -6250 16600 -5350 16700
rect -4850 16650 -4700 16750
rect -4300 16800 -3500 16950
rect -4300 16700 -3450 16800
rect -4900 16600 -4700 16650
rect -8000 16500 -6800 16600
rect -6300 16500 -5400 16600
rect -4900 16550 -4650 16600
rect -8000 16400 -6850 16500
rect -6350 16450 -5400 16500
rect -4950 16450 -4650 16550
rect -4250 16450 -3450 16700
rect -6350 16400 -5450 16450
rect -8000 16300 -6900 16400
rect -6400 16350 -5450 16400
rect -5000 16350 -4650 16450
rect -6400 16300 -5500 16350
rect -8000 16200 -6950 16300
rect -6450 16250 -5500 16300
rect -5050 16250 -4600 16350
rect -8000 16100 -7000 16200
rect -6450 16150 -5550 16250
rect -8000 16050 -7050 16100
rect -6500 16050 -5600 16150
rect -5100 16100 -4600 16250
rect -4200 16300 -3450 16450
rect -4200 16200 -3500 16300
rect -7950 16000 -7050 16050
rect -7950 15900 -7100 16000
rect -6550 15950 -6100 16050
rect -6000 16000 -5650 16050
rect -5150 16000 -4550 16100
rect -5900 15950 -5650 16000
rect -6600 15900 -6100 15950
rect -5750 15900 -5700 15950
rect -5200 15900 -4550 16000
rect -4150 16000 -3500 16200
rect -4150 15950 -3550 16000
rect -7950 15850 -7150 15900
rect -6600 15850 -6150 15900
rect -5250 15850 -4550 15900
rect -7900 15750 -7150 15850
rect -5300 15750 -4500 15850
rect -4100 15800 -3550 15950
rect -4100 15750 -3600 15800
rect -7900 15700 -7200 15750
rect -5200 15700 -4500 15750
rect -7850 15650 -7200 15700
rect -5050 15650 -4500 15700
rect -7850 15550 -7250 15650
rect -4900 15600 -4500 15650
rect -4050 15650 -3600 15750
rect -4750 15550 -4450 15600
rect -7800 15450 -7300 15550
rect -4950 15500 -4450 15550
rect -4050 15550 -3650 15650
rect -4050 15500 -3700 15550
rect -5100 15450 -4450 15500
rect -7750 15400 -7350 15450
rect -5300 15400 -4450 15450
rect -7750 15350 -7400 15400
rect -5500 15350 -4450 15400
rect -4000 15450 -3700 15500
rect -4000 15350 -3750 15450
rect -7700 15300 -6400 15350
rect -5650 15300 -4400 15350
rect -7650 15250 -6400 15300
rect -5850 15250 -4400 15300
rect -4000 15250 -3800 15350
rect -7650 15200 -6450 15250
rect -6050 15200 -4400 15250
rect -7600 15150 -6500 15200
rect -6200 15150 -5650 15200
rect -5550 15150 -4400 15200
rect -3950 15150 -3850 15250
rect -7550 15100 -6500 15150
rect -6400 15100 -5750 15150
rect -7550 15050 -5900 15100
rect -5600 15050 -4350 15150
rect -7500 15000 -6000 15050
rect -7450 14950 -6100 15000
rect -5650 14950 -4350 15050
rect -7400 14900 -6150 14950
rect -5700 14900 -4350 14950
rect -7350 14850 -6200 14900
rect -5700 14850 -4300 14900
rect -7300 14800 -6200 14850
rect -7250 14750 -6250 14800
rect -5750 14750 -4300 14850
rect -7200 14700 -6250 14750
rect -7150 14650 -6300 14700
rect -5800 14650 -4300 14750
rect -7100 14600 -6300 14650
rect -5850 14600 -4400 14650
rect -7050 14550 -6350 14600
rect -5850 14550 -4450 14600
rect -6950 14500 -6350 14550
rect -5900 14500 -4550 14550
rect -6900 14450 -6400 14500
rect -5900 14450 -4600 14500
rect -6800 14400 -6400 14450
rect -5950 14400 -4700 14450
rect -6700 14350 -6450 14400
rect -5950 14350 -4800 14400
rect -6600 14300 -6450 14350
rect -6000 14300 -4900 14350
rect -6000 14250 -5050 14300
rect -6050 14200 -5200 14250
rect -6050 14150 -5450 14200
rect -8700 13550 -8600 13600
rect -9150 13500 -8600 13550
rect -7500 13500 -7400 13600
rect -9000 13400 -8900 13500
rect -8750 13461 -8600 13500
rect -8750 13450 -8582 13461
rect -7550 13450 -7400 13500
rect -5500 13450 -5350 13550
rect -5200 13500 -5050 13550
rect -8750 13400 -8650 13450
rect -8613 13437 -8450 13450
rect -8600 13411 -8450 13437
rect -8300 13412 -8100 13450
rect -8613 13400 -8450 13411
rect -8314 13400 -8100 13412
rect -7950 13400 -7650 13450
rect -9050 13200 -8950 13400
rect -8750 13384 -8584 13400
rect -8750 13350 -8600 13384
rect -8750 13250 -8650 13350
rect -8550 13250 -8450 13400
rect -8350 13384 -8289 13400
rect -8350 13350 -8300 13384
rect -8150 13300 -8050 13400
rect -7950 13300 -7850 13400
rect -8350 13250 -8050 13300
rect -8800 13200 -8650 13250
rect -9100 13100 -9000 13200
rect -8800 13100 -8700 13200
rect -8600 13100 -8500 13250
rect -8400 13150 -8300 13250
rect -8150 13200 -8050 13250
rect -8000 13250 -7850 13300
rect -7750 13250 -7650 13400
rect -7550 13350 -7450 13450
rect -7350 13400 -7250 13450
rect -7400 13350 -7300 13400
rect -7550 13250 -7350 13350
rect -6950 13300 -6850 13450
rect -6700 13400 -6600 13450
rect -6500 13400 -6300 13450
rect -6750 13300 -6650 13400
rect -6550 13350 -6450 13400
rect -8200 13150 -8100 13200
rect -8400 13100 -8100 13150
rect -8000 13100 -7900 13250
rect -7800 13100 -7700 13250
rect -7600 13200 -7350 13250
rect -6900 13200 -6700 13300
rect -7600 13100 -7500 13200
rect -7400 13150 -7300 13200
rect -7400 13100 -7250 13150
rect -6900 13100 -6750 13200
rect -6600 13150 -6500 13350
rect -6350 13200 -6250 13400
rect -6150 13300 -6050 13450
rect -5950 13300 -5850 13450
rect -6400 13150 -6300 13200
rect -6200 13150 -6100 13300
rect -6000 13250 -5850 13300
rect -6000 13150 -5900 13250
rect -5550 13200 -5450 13450
rect -5400 13300 -5350 13450
rect -5250 13450 -5050 13500
rect -4500 13450 -4400 13500
rect -4200 13450 -4100 13500
rect -5250 13400 -5100 13450
rect -4900 13420 -4700 13450
rect -4920 13400 -4700 13420
rect -4550 13400 -4300 13450
rect -4250 13400 -4000 13450
rect -3750 13400 -3650 13550
rect -3450 13500 -3300 13550
rect -3450 13450 -3350 13500
rect -3500 13417 -3350 13450
rect -3500 13400 -3369 13417
rect -3300 13400 -3100 13450
rect -2950 13400 -2650 13450
rect -5300 13350 -5100 13400
rect -4950 13381 -4884 13400
rect -4950 13350 -4900 13381
rect -5300 13300 -5250 13350
rect -5400 13250 -5250 13300
rect -5400 13200 -5300 13250
rect -5200 13200 -5100 13350
rect -4750 13300 -4650 13400
rect -4500 13350 -4400 13400
rect -4200 13350 -4100 13400
rect -4950 13250 -4650 13300
rect -6550 13100 -6350 13150
rect -6200 13100 -5900 13150
rect -5600 13100 -5500 13200
rect -5250 13100 -5150 13200
rect -5000 13150 -4900 13250
rect -4750 13200 -4650 13250
rect -4550 13300 -4400 13350
rect -4250 13300 -4100 13350
rect -4800 13150 -4700 13200
rect -5000 13100 -4700 13150
rect -4550 13150 -4450 13300
rect -4250 13150 -4150 13300
rect -3700 13250 -3600 13400
rect -3500 13366 -3400 13400
rect -3326 13384 -3250 13400
rect -3500 13350 -3423 13366
rect -3350 13350 -3250 13384
rect -3550 13250 -3450 13350
rect -3382 13330 -3300 13350
rect -3400 13300 -3300 13330
rect -3150 13300 -3050 13400
rect -2950 13300 -2850 13400
rect -3400 13250 -3050 13300
rect -3000 13250 -2850 13300
rect -2750 13250 -2650 13400
rect -2550 13400 -2250 13450
rect -2550 13300 -2450 13400
rect -2600 13250 -2450 13300
rect -2350 13250 -2250 13400
rect -3700 13150 -3500 13250
rect -3400 13150 -3300 13250
rect -3150 13170 -3100 13200
rect -3176 13150 -3100 13170
rect -4550 13100 -4350 13150
rect -4250 13100 -4050 13150
rect -3700 13100 -3550 13150
rect -3350 13127 -3125 13150
rect -3350 13100 -3150 13127
rect -3000 13100 -2900 13250
rect -2800 13100 -2700 13250
rect -2600 13100 -2500 13250
rect -2400 13100 -2300 13250
rect -6900 13000 -6800 13100
rect -7000 12950 -6850 13000
rect -7450 12600 -7350 12800
rect -7150 12750 -7050 12800
rect -6650 12750 -6550 12850
rect -6200 12769 -6000 12800
rect -6221 12750 -6000 12769
rect -5800 12750 -5700 12850
rect -5000 12750 -4900 12850
rect -4000 12750 -3900 12850
rect -7500 12400 -7400 12600
rect -7200 12500 -7100 12750
rect -6300 12728 -6178 12750
rect -7000 12650 -6750 12700
rect -7000 12550 -6900 12650
rect -6700 12550 -6600 12700
rect -6300 12650 -6200 12728
rect -6050 12700 -6000 12750
rect -5850 12726 -5700 12750
rect -5850 12700 -5677 12726
rect -5050 12700 -4900 12750
rect -4050 12700 -3900 12750
rect -5850 12650 -5750 12700
rect -5717 12667 -5550 12700
rect -5400 12672 -5200 12700
rect -5720 12650 -5550 12667
rect -5419 12650 -5200 12672
rect -6300 12600 -6150 12650
rect -5850 12622 -5679 12650
rect -5850 12600 -5700 12622
rect -6250 12550 -6000 12600
rect -7050 12500 -6900 12550
rect -6750 12500 -6600 12550
rect -6150 12500 -6000 12550
rect -5850 12500 -5750 12600
rect -5650 12500 -5550 12650
rect -5450 12634 -5381 12650
rect -5450 12600 -5400 12634
rect -5250 12550 -5150 12650
rect -5450 12500 -5150 12550
rect -5050 12600 -4950 12700
rect -4850 12650 -4750 12700
rect -4600 12650 -4400 12700
rect -4200 12650 -3950 12700
rect -4900 12600 -4800 12650
rect -4650 12600 -4550 12650
rect -5050 12500 -4850 12600
rect -7250 12400 -7150 12500
rect -7450 12350 -7200 12400
rect -7050 12350 -6950 12500
rect -6750 12350 -6650 12500
rect -6350 12400 -6300 12450
rect -6100 12400 -6000 12500
rect -5900 12450 -5750 12500
rect -6350 12350 -6050 12400
rect -5900 12350 -5800 12450
rect -5700 12350 -5600 12500
rect -5500 12400 -5400 12500
rect -5250 12450 -5150 12500
rect -5100 12450 -4850 12500
rect -4700 12550 -4600 12600
rect -4450 12550 -4350 12650
rect -4250 12600 -4150 12650
rect -4700 12500 -4350 12550
rect -5300 12400 -5200 12450
rect -5500 12350 -5200 12400
rect -5100 12350 -5000 12450
rect -4900 12400 -4800 12450
rect -4700 12400 -4600 12500
rect -4450 12419 -4400 12450
rect -4467 12400 -4400 12419
rect -4300 12400 -4200 12600
rect -4050 12500 -3950 12650
rect -4100 12450 -3950 12500
rect -4100 12400 -4000 12450
rect -4900 12350 -4750 12400
rect -4650 12381 -4432 12400
rect -4650 12350 -4450 12381
rect -4250 12350 -4000 12400
rect -8250 12050 -8000 12100
rect -7750 12050 -7650 12150
rect -6050 12062 -5850 12100
rect -6064 12050 -5850 12062
rect -4950 12050 -4850 12150
rect -4000 12050 -3900 12150
rect -3150 12050 -3050 12150
rect -8250 12000 -8150 12050
rect -8050 12000 -7950 12050
rect -6150 12030 -6029 12050
rect -8300 11750 -8200 12000
rect -8000 11800 -7900 12000
rect -7800 11850 -7700 12000
rect -7550 11950 -7350 12000
rect -7150 11950 -6850 12000
rect -6700 11950 -6500 12000
rect -6150 11950 -6050 12030
rect -5900 12000 -5850 12050
rect -5250 12000 -5150 12050
rect -4050 12017 -3900 12050
rect -4050 12000 -3880 12017
rect -3200 12000 -3050 12050
rect -5650 11971 -5450 12000
rect -5669 11950 -5450 11971
rect -5300 11950 -5050 12000
rect -7600 11900 -7500 11950
rect -7850 11800 -7700 11850
rect -7650 11850 -7550 11900
rect -7400 11850 -7300 11950
rect -7200 11900 -7100 11950
rect -7650 11800 -7300 11850
rect -8050 11750 -7950 11800
rect -8350 11700 -8250 11750
rect -8100 11700 -7950 11750
rect -8350 11650 -8050 11700
rect -7850 11650 -7750 11800
rect -7650 11700 -7550 11800
rect -7400 11721 -7350 11750
rect -7421 11700 -7350 11721
rect -7250 11700 -7150 11900
rect -7000 11850 -6850 11950
rect -6750 11900 -6650 11950
rect -7000 11750 -6900 11850
rect -7050 11716 -6900 11750
rect -7061 11700 -6900 11716
rect -6800 11700 -6700 11900
rect -6550 11750 -6450 11950
rect -6150 11900 -6000 11950
rect -5700 11933 -5629 11950
rect -5700 11900 -5650 11933
rect -6100 11850 -5850 11900
rect -5500 11850 -5400 11950
rect -5250 11900 -5150 11950
rect -6000 11800 -5850 11850
rect -5700 11800 -5400 11850
rect -6600 11700 -6500 11750
rect -6200 11700 -6150 11750
rect -5950 11700 -5850 11800
rect -5750 11700 -5650 11800
rect -5500 11750 -5400 11800
rect -5300 11850 -5150 11900
rect -5000 11850 -4900 12000
rect -4800 11950 -4500 12000
rect -4400 11971 -4200 12000
rect -4414 11950 -4200 11971
rect -4050 11950 -3950 12000
rect -3918 11986 -3750 12000
rect -3899 11967 -3750 11986
rect -3550 11974 -3350 12000
rect -3920 11950 -3750 11967
rect -3566 11950 -3350 11974
rect -4650 11900 -4500 11950
rect -4450 11928 -4378 11950
rect -4450 11900 -4400 11928
rect -4700 11850 -4550 11900
rect -4250 11850 -4150 11950
rect -5550 11700 -5450 11750
rect -7600 11678 -7380 11700
rect -7200 11690 -7036 11700
rect -7600 11650 -7400 11678
rect -7200 11668 -7050 11690
rect -7200 11650 -7026 11668
rect -7000 11650 -6900 11700
rect -6750 11650 -6550 11700
rect -6200 11650 -5900 11700
rect -5750 11650 -5450 11700
rect -5300 11700 -5200 11850
rect -5050 11800 -4900 11850
rect -4750 11800 -4600 11850
rect -4450 11800 -4150 11850
rect -4050 11936 -3882 11950
rect -4050 11900 -3900 11936
rect -4050 11800 -3950 11900
rect -5300 11650 -5100 11700
rect -5050 11650 -4950 11800
rect -4800 11750 -4650 11800
rect -4850 11700 -4700 11750
rect -4500 11700 -4400 11800
rect -4250 11750 -4150 11800
rect -4300 11700 -4200 11750
rect -4850 11650 -4550 11700
rect -4500 11650 -4200 11700
rect -4100 11700 -3950 11800
rect -3800 11750 -3700 11950
rect -3600 11931 -3528 11950
rect -3600 11900 -3550 11931
rect -3400 11850 -3300 11950
rect -3600 11800 -3300 11850
rect -3200 11800 -3100 12000
rect -3850 11700 -3750 11750
rect -3650 11700 -3550 11800
rect -3400 11750 -3300 11800
rect -3250 11750 -3100 11800
rect -3450 11700 -3350 11750
rect -4100 11650 -3800 11700
rect -3650 11650 -3350 11700
rect -3250 11650 -3150 11750
rect -7066 11630 -6950 11650
rect -7250 11550 -7200 11600
rect -7050 11550 -6950 11630
rect -7250 11500 -7000 11550
rect -8050 11350 -7950 11400
rect -8500 11300 -7950 11350
rect -7100 11300 -6650 11350
rect -8350 11200 -8250 11300
rect -8400 11000 -8300 11200
rect -8100 11100 -8000 11250
rect -7900 11200 -7600 11250
rect -7900 11100 -7800 11200
rect -8150 11050 -8000 11100
rect -7950 11050 -7800 11100
rect -7700 11050 -7600 11200
rect -7500 11100 -7400 11250
rect -7250 11200 -7150 11250
rect -6950 11200 -6850 11300
rect -4700 11250 -4600 11300
rect -6700 11220 -6500 11250
rect -6712 11200 -6500 11220
rect -6350 11200 -6100 11250
rect -5900 11200 -5700 11250
rect -5500 11200 -5300 11250
rect -7300 11100 -7200 11200
rect -8450 10900 -8350 11000
rect -8150 10900 -8050 11050
rect -7950 10900 -7850 11050
rect -7750 10900 -7650 11050
rect -7450 11000 -7250 11100
rect -7000 11000 -6900 11200
rect -6750 11177 -6677 11200
rect -6750 11150 -6700 11177
rect -6550 11100 -6450 11200
rect -6350 11150 -6250 11200
rect -6750 11050 -6450 11100
rect -7450 10900 -7300 11000
rect -7050 10900 -6950 11000
rect -6800 10950 -6700 11050
rect -6550 11000 -6450 11050
rect -6400 11100 -6250 11150
rect -6600 10950 -6500 11000
rect -6800 10900 -6500 10950
rect -6400 10950 -6300 11100
rect -6150 11000 -6050 11200
rect -5950 11150 -5850 11200
rect -6000 11100 -5900 11150
rect -5750 11100 -5650 11200
rect -5550 11150 -5450 11200
rect -6000 11050 -5650 11100
rect -6200 10950 -6100 11000
rect -6000 10950 -5900 11050
rect -5750 10974 -5700 11000
rect -5771 10950 -5700 10974
rect -5600 10950 -5500 11150
rect -5350 11000 -5250 11200
rect -5150 11100 -5050 11250
rect -4950 11100 -4850 11250
rect -4750 11200 -4500 11250
rect -4150 11214 -3950 11250
rect -4150 11200 -3935 11214
rect -3800 11200 -3600 11250
rect -3450 11200 -2900 11250
rect -4700 11150 -4600 11200
rect -4200 11150 -4100 11200
rect -3968 11179 -3900 11200
rect -3950 11169 -3900 11179
rect -3950 11150 -3918 11169
rect -3850 11150 -3750 11200
rect -5400 10950 -5300 11000
rect -5200 10950 -5100 11100
rect -5000 11050 -4850 11100
rect -4750 11100 -4600 11150
rect -5000 10950 -4900 11050
rect -6400 10900 -6150 10950
rect -5950 10931 -5733 10950
rect -5950 10900 -5750 10931
rect -5550 10900 -5350 10950
rect -5200 10900 -4900 10950
rect -4750 10950 -4650 11100
rect -4750 10900 -4550 10950
rect -4450 10900 -4350 11000
rect -4250 10950 -4150 11150
rect -3882 11136 -3800 11150
rect -4000 10972 -3950 11000
rect -4022 10950 -3950 10972
rect -3900 10950 -3800 11136
rect -3650 11000 -3550 11200
rect -3450 11100 -3350 11200
rect -3500 11050 -3350 11100
rect -3200 11050 -3100 11200
rect -3000 11050 -2900 11200
rect -3700 10950 -3600 11000
rect -4200 10936 -3984 10950
rect -4200 10900 -4000 10936
rect -3850 10900 -3650 10950
rect -3500 10900 -3400 11050
rect -3250 11000 -3100 11050
rect -3250 10900 -3150 11000
rect -3050 10900 -2950 11050
rect -7450 10800 -7350 10900
rect -6450 10850 -6300 10900
rect -7550 10750 -7400 10800
rect -6450 10750 -6350 10850
rect -9000 10600 -8600 10650
rect -6200 10600 -6050 10650
rect -5800 10620 -5600 10650
rect -5824 10600 -5600 10620
rect -8750 10550 -8600 10600
rect -7200 10550 -7100 10600
rect -6250 10550 -6050 10600
rect -8800 10500 -8650 10550
rect -8500 10500 -8300 10550
rect -8150 10500 -7900 10550
rect -7800 10500 -7600 10550
rect -7250 10500 -7000 10550
rect -6900 10500 -6700 10550
rect -6250 10500 -6200 10550
rect -8850 10450 -8700 10500
rect -8550 10450 -8450 10500
rect -8900 10400 -8750 10450
rect -8600 10400 -8500 10450
rect -8350 10400 -8250 10500
rect -8150 10400 -8050 10500
rect -7850 10450 -7750 10500
rect -8950 10350 -8800 10400
rect -8600 10350 -8250 10400
rect -8200 10350 -8050 10400
rect -9000 10300 -8850 10350
rect -9050 10250 -8900 10300
rect -8600 10250 -8500 10350
rect -8350 10268 -8300 10300
rect -8365 10250 -8300 10268
rect -9050 10200 -8650 10250
rect -8550 10235 -8329 10250
rect -8550 10200 -8350 10235
rect -8200 10200 -8100 10350
rect -7900 10250 -7800 10450
rect -7650 10300 -7550 10500
rect -7200 10450 -7100 10500
rect -6950 10450 -6850 10500
rect -7250 10400 -7100 10450
rect -7700 10250 -7600 10300
rect -7250 10250 -7150 10400
rect -7000 10250 -6900 10450
rect -6750 10300 -6650 10500
rect -6300 10400 -6200 10500
rect -6350 10350 -6250 10400
rect -6150 10350 -6050 10550
rect -5900 10582 -5783 10600
rect -5900 10500 -5800 10582
rect -5650 10550 -5600 10600
rect -5400 10550 -5300 10650
rect -5150 10600 -4900 10650
rect -4500 10600 -4250 10650
rect -5200 10550 -5100 10600
rect -4950 10550 -4900 10600
rect -4550 10550 -4450 10600
rect -4300 10550 -4250 10600
rect -5900 10450 -5750 10500
rect -5850 10400 -5600 10450
rect -5750 10350 -5600 10400
rect -6400 10300 -6000 10350
rect -6800 10250 -6700 10300
rect -6400 10250 -6300 10300
rect -7850 10200 -7650 10250
rect -7250 10200 -7050 10250
rect -6950 10200 -6750 10250
rect -6450 10200 -6300 10250
rect -6100 10200 -6000 10300
rect -5950 10250 -5900 10300
rect -5700 10250 -5600 10350
rect -5450 10300 -5350 10550
rect -5250 10500 -5150 10550
rect -4600 10500 -4500 10550
rect -4100 10500 -3900 10550
rect -5300 10300 -5200 10500
rect -4650 10300 -4550 10500
rect -4150 10450 -4050 10500
rect -5950 10200 -5650 10250
rect -5500 10200 -5400 10300
rect -5250 10250 -5150 10300
rect -5000 10250 -4950 10300
rect -4600 10250 -4500 10300
rect -4350 10250 -4300 10300
rect -4200 10250 -4100 10450
rect -3950 10300 -3850 10500
rect -3750 10400 -3650 10550
rect -3550 10400 -3450 10550
rect -3350 10500 -3100 10550
rect -3000 10500 -2800 10550
rect -2650 10500 -2450 10550
rect -3350 10400 -3250 10500
rect -4000 10250 -3900 10300
rect -3800 10250 -3700 10400
rect -3600 10350 -3450 10400
rect -3400 10350 -3250 10400
rect -3050 10450 -2950 10500
rect -2850 10450 -2800 10500
rect -2700 10450 -2600 10500
rect -3050 10400 -2900 10450
rect -2750 10400 -2650 10450
rect -2500 10400 -2400 10500
rect -3050 10350 -2800 10400
rect -3600 10250 -3500 10350
rect -5200 10200 -4950 10250
rect -4550 10200 -4300 10250
rect -4150 10200 -3950 10250
rect -3800 10200 -3500 10250
rect -3400 10200 -3300 10350
rect -2950 10300 -2800 10350
rect -3100 10275 -3050 10300
rect -3100 10250 -3034 10275
rect -2900 10250 -2800 10300
rect -2750 10350 -2400 10400
rect -2750 10250 -2650 10350
rect -2500 10275 -2450 10300
rect -2521 10250 -2450 10275
rect -3075 10232 -2850 10250
rect -3050 10200 -2850 10232
rect -2700 10232 -2480 10250
rect -2700 10200 -2500 10232
rect -8550 9900 -8400 9950
rect -8600 9850 -8400 9900
rect -6900 9900 -6650 9950
rect -4150 9919 -3950 9950
rect -4171 9900 -3950 9919
rect -3750 9900 -3550 9950
rect -3350 9921 -3150 9950
rect -3374 9900 -3150 9921
rect -2850 9900 -2700 9950
rect -6900 9850 -6800 9900
rect -6700 9850 -6600 9900
rect -4250 9881 -4125 9900
rect -4250 9850 -4150 9881
rect -8600 9800 -8550 9850
rect -8650 9700 -8550 9800
rect -8700 9650 -8600 9700
rect -8500 9650 -8400 9850
rect -8250 9800 -8000 9850
rect -7900 9800 -7700 9850
rect -7550 9800 -7250 9850
rect -8250 9700 -8150 9800
rect -7950 9750 -7850 9800
rect -8300 9650 -8150 9700
rect -8750 9600 -8350 9650
rect -8750 9550 -8650 9600
rect -8800 9500 -8650 9550
rect -8450 9500 -8350 9600
rect -8300 9500 -8200 9650
rect -8000 9550 -7900 9750
rect -7750 9600 -7650 9800
rect -7550 9700 -7450 9800
rect -7600 9650 -7450 9700
rect -7350 9650 -7250 9800
rect -7800 9550 -7700 9600
rect -7950 9500 -7750 9550
rect -7600 9500 -7500 9650
rect -7400 9500 -7300 9650
rect -6950 9600 -6850 9850
rect -6650 9650 -6550 9850
rect -6400 9800 -6200 9850
rect -6050 9800 -5750 9850
rect -6450 9750 -6350 9800
rect -6500 9700 -6400 9750
rect -6250 9700 -6150 9800
rect -6050 9700 -5950 9800
rect -6500 9650 -6150 9700
rect -6100 9650 -5950 9700
rect -5850 9650 -5750 9800
rect -5650 9800 -5350 9850
rect -5200 9800 -5000 9850
rect -4850 9800 -4550 9850
rect -5650 9700 -5550 9800
rect -5700 9650 -5550 9700
rect -5450 9650 -5350 9800
rect -5250 9750 -5150 9800
rect -5300 9700 -5200 9750
rect -5050 9700 -4950 9800
rect -4850 9700 -4750 9800
rect -5300 9650 -4950 9700
rect -4900 9650 -4750 9700
rect -4650 9650 -4550 9800
rect -4000 9750 -3900 9900
rect -3800 9800 -3700 9900
rect -4050 9700 -3950 9750
rect -4150 9650 -4000 9700
rect -6700 9600 -6600 9650
rect -7000 9550 -6900 9600
rect -6750 9550 -6600 9600
rect -6500 9550 -6400 9650
rect -6250 9572 -6200 9600
rect -6272 9550 -6200 9572
rect -7000 9500 -6700 9550
rect -6450 9526 -6231 9550
rect -6450 9500 -6250 9526
rect -6100 9500 -6000 9650
rect -5900 9500 -5800 9650
rect -5700 9500 -5600 9650
rect -5500 9500 -5400 9650
rect -5300 9550 -5200 9650
rect -5050 9574 -5000 9600
rect -5067 9550 -5000 9574
rect -5250 9531 -5029 9550
rect -5250 9500 -5050 9531
rect -4900 9500 -4800 9650
rect -4700 9500 -4600 9650
rect -4200 9600 -4100 9650
rect -4300 9550 -4150 9600
rect -3850 9550 -3750 9800
rect -3600 9650 -3500 9900
rect -3450 9881 -3328 9900
rect -3450 9850 -3350 9881
rect -3200 9750 -3100 9900
rect -2900 9850 -2700 9900
rect -2900 9820 -2750 9850
rect -2920 9800 -2750 9820
rect -2950 9779 -2882 9800
rect -2950 9750 -2900 9779
rect -3250 9700 -3150 9750
rect -3000 9700 -2900 9750
rect -3350 9650 -3200 9700
rect -3050 9650 -2950 9700
rect -2850 9650 -2750 9800
tri -1250 9650 -1100 9800 se
rect -1100 9650 -100 9800
rect -3650 9550 -3550 9650
rect -3400 9600 -3300 9650
rect -3050 9600 -2700 9650
tri -1300 9600 -1250 9650 se
rect -1250 9600 -100 9650
rect -3500 9550 -3350 9600
rect -4300 9500 -3950 9550
rect -3800 9500 -3600 9550
rect -3500 9500 -3150 9550
rect -2900 9500 -2800 9600
tri -1400 9500 -1300 9600 se
rect -1300 9500 -100 9600
tri -1600 9300 -1400 9500 se
rect -1400 9300 -100 9500
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -4207 4950 -3500 5657 se
tri -3500 4950 -2793 5657 sw
tri -4207 4243 -3500 4950 ne
tri -3500 4243 -2793 4950 nw
rect 0 500 200 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal3 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -4207 6450 -3500 7157 se
tri -3500 6450 -2793 7157 sw
tri -4207 5743 -3500 6450 ne
tri -3500 5743 -2793 6450 nw
rect 300 500 500 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal4 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
tri -4207 7950 -3500 8657 se
tri -3500 7950 -2793 8657 sw
tri -4207 7243 -3500 7950 ne
tri -3500 7243 -2793 7950 nw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
rect 600 500 800 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< end >>

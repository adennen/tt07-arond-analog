magic
tech sky130A
timestamp 1717261812
<< metal1 >>
rect -300 500 -100 700
tri -200 300 -100 400 se
tri -100 300 0 400 sw
rect 500 300 800 400
tri 800 300 900 400 sw
tri -300 200 -200 300 se
tri -200 200 -100 300 nw
tri -100 200 0 300 ne
tri 0 200 100 300 sw
tri -500 0 -300 200 se
tri -300 100 -200 200 nw
tri 0 100 100 200 ne
tri 100 100 200 200 sw
rect 100 0 200 100
tri 200 0 300 100 sw
rect -500 -100 300 0
rect -500 -200 -300 -100
rect 100 -200 300 -100
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal2 >>
rect 0 500 200 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal3 >>
rect 300 500 500 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal4 >>
rect 600 500 800 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< end >>

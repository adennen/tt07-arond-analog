magic
tech sky130A
timestamp 1717265593
<< metal1 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -1100 5300 -100 6300 se
rect -100 5300 900 6300
tri -1600 4800 -1100 5300 se
tri -1100 4800 -600 5300 nw
tri -2100 4300 -1600 4800 se
tri -1600 4300 -1100 4800 nw
tri -2100 4157 -1957 4300 ne
rect -1957 4157 -1600 4300
tri -4207 3450 -3500 4157 se
tri -3500 3450 -2793 4157 sw
tri -1957 3800 -1600 4157 ne
tri -1600 3800 -1100 4300 sw
tri -4207 2743 -3500 3450 ne
tri -3500 2743 -2793 3450 nw
tri -1600 3300 -1100 3800 ne
tri -1100 3300 -600 3800 sw
rect -100 3300 400 5300
tri -1100 2743 -543 3300 ne
rect -543 2743 900 3300
tri -543 2300 -100 2743 ne
rect -100 2300 900 2743
rect -300 500 -100 700
tri -200 300 -100 400 se
tri -100 300 0 400 sw
rect 500 300 800 400
tri 800 300 900 400 sw
tri -300 200 -200 300 se
tri -200 200 -100 300 nw
tri -100 200 0 300 ne
tri 0 200 100 300 sw
tri -500 0 -300 200 se
tri -300 100 -200 200 nw
tri 0 100 100 200 ne
tri 100 100 200 200 sw
rect 100 0 200 100
tri 200 0 300 100 sw
rect -500 -100 300 0
rect -500 -200 -300 -100
rect 100 -200 300 -100
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal2 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -4207 4950 -3500 5657 se
tri -3500 4950 -2793 5657 sw
tri -4207 4243 -3500 4950 ne
tri -3500 4243 -2793 4950 nw
rect 0 500 200 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal3 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
tri -4207 6450 -3500 7157 se
tri -3500 6450 -2793 7157 sw
tri -4207 5743 -3500 6450 ne
tri -3500 5743 -2793 6450 nw
rect 300 500 500 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< metal4 >>
tri -1600 9300 -1100 9800 se
rect -1100 9300 -100 9800
tri -100 9300 400 9800 sw
tri -2100 8800 -1600 9300 se
tri -1600 8800 -1100 9300 nw
tri -100 8800 400 9300 ne
tri 400 8800 900 9300 sw
tri -4207 7950 -3500 8657 se
tri -3500 7950 -2793 8657 sw
tri -4207 7243 -3500 7950 ne
tri -3500 7243 -2793 7950 nw
rect -2100 7800 -1600 8800
rect 400 7800 900 8800
rect -2100 7300 900 7800
rect 600 500 800 700
rect 500 300 800 400
tri 800 300 900 400 sw
rect 500 -100 600 300
tri 800 200 900 300 ne
tri 900 200 1000 300 sw
rect 900 0 1000 200
tri 800 -100 900 0 se
tri 900 -100 1000 0 nw
rect 500 -200 800 -100
tri 800 -200 900 -100 nw
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1717269404
<< metal1 >>
rect 25940 3392 26240 3398
rect 26240 3092 27198 3392
rect 25940 3086 26240 3092
rect 26866 2068 27046 2258
rect 31282 2074 31462 2266
rect 26860 1888 26866 2068
rect 27046 1888 27052 2068
rect 31276 1894 31282 2074
rect 31462 1894 31468 2074
rect 25938 1322 26238 1328
rect 26238 1022 27132 1322
rect 25938 1016 26238 1022
<< via1 >>
rect 25940 3092 26240 3392
rect 26866 1888 27046 2068
rect 31282 1894 31462 2074
rect 25938 1022 26238 1322
<< metal2 >>
rect 25347 3392 25637 3396
rect 25342 3387 25940 3392
rect 25342 3097 25347 3387
rect 25637 3097 25940 3387
rect 25342 3092 25940 3097
rect 26240 3092 26246 3392
rect 25347 3088 25637 3092
rect 31282 2074 31462 2080
rect 26866 2068 27046 2074
rect 26866 1879 27046 1888
rect 26862 1709 26871 1879
rect 27041 1709 27050 1879
rect 31282 1873 31462 1894
rect 26866 1704 27046 1709
rect 31278 1703 31287 1873
rect 31457 1703 31466 1873
rect 31282 1698 31462 1703
rect 25341 1322 25631 1326
rect 25336 1317 25938 1322
rect 25336 1027 25341 1317
rect 25631 1027 25938 1317
rect 25336 1022 25938 1027
rect 26238 1022 26244 1322
rect 25341 1018 25631 1022
<< via2 >>
rect 25347 3097 25637 3387
rect 26871 1709 27041 1879
rect 31287 1703 31457 1873
rect 25341 1027 25631 1317
<< metal3 >>
rect 7683 3392 7981 3397
rect 24697 3392 24995 3397
rect 7682 3391 11462 3392
rect 7682 3093 7683 3391
rect 7981 3093 11462 3391
rect 7682 3092 11462 3093
rect 11762 3092 11768 3392
rect 24696 3391 25642 3392
rect 24696 3093 24697 3391
rect 24995 3387 25642 3391
rect 24995 3097 25347 3387
rect 25637 3097 25642 3387
rect 24995 3093 25642 3097
rect 24696 3092 25642 3093
rect 7683 3087 7981 3092
rect 24697 3087 24995 3092
rect 26866 1879 27046 1884
rect 26866 1709 26871 1879
rect 27041 1709 27046 1879
rect 31282 1873 31462 1878
rect 31282 1721 31287 1873
rect 31457 1721 31462 1873
rect 26866 1707 27046 1709
rect 26861 1529 26867 1707
rect 27045 1529 27051 1707
rect 31277 1543 31283 1721
rect 31461 1543 31467 1721
rect 31282 1542 31462 1543
rect 26866 1528 27046 1529
rect 24685 1322 24983 1327
rect 24684 1321 25636 1322
rect 24684 1023 24685 1321
rect 24983 1317 25636 1321
rect 24983 1027 25341 1317
rect 25631 1027 25636 1317
rect 24983 1023 25636 1027
rect 24684 1022 25636 1023
rect 24685 1017 24983 1022
<< via3 >>
rect 7683 3093 7981 3391
rect 11462 3092 11762 3392
rect 24697 3093 24995 3391
rect 26867 1529 27045 1707
rect 31283 1703 31287 1721
rect 31287 1703 31457 1721
rect 31457 1703 31461 1721
rect 31283 1543 31461 1703
rect 24685 1023 24983 1321
<< metal4 >>
rect 798 44742 858 45152
rect 1534 44742 1594 45152
rect 2270 44742 2330 45152
rect 3006 44742 3066 45152
rect 3742 44742 3802 45152
rect 4478 44742 4538 45152
rect 5214 44742 5274 45152
rect 5950 44742 6010 45152
rect 6686 44742 6746 45152
rect 7422 44742 7482 45152
rect 8158 44742 8218 45152
rect 8894 44742 8954 45152
rect 9630 44742 9690 45152
rect 10366 44742 10426 45152
rect 11102 44742 11162 45152
rect 11838 44742 11898 45152
rect 12574 44742 12634 45152
rect 13310 44742 13370 45152
rect 14046 44742 14106 45152
rect 14782 44742 14842 45152
rect 15518 44742 15578 45152
rect 16254 44742 16314 45152
rect 16990 44742 17050 45152
rect 17726 44742 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 400 44526 18094 44742
rect 9838 44152 10054 44526
rect 200 3392 500 44152
rect 200 3391 7982 3392
rect 200 3093 7683 3391
rect 7981 3093 7982 3391
rect 200 3092 7982 3093
rect 200 1000 500 3092
rect 9800 1322 10100 44152
rect 11461 3392 11763 3393
rect 11461 3092 11462 3392
rect 11762 3391 24996 3392
rect 11762 3093 24697 3391
rect 24995 3093 24996 3391
rect 11762 3092 24996 3093
rect 11461 3091 11763 3092
rect 31282 1721 31462 1722
rect 26866 1707 27046 1708
rect 26866 1529 26867 1707
rect 27045 1529 27046 1707
rect 9800 1321 24984 1322
rect 9800 1023 24685 1321
rect 24983 1023 24984 1321
rect 9800 1022 24984 1023
rect 9800 1000 10100 1022
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 1529
rect 31282 1543 31283 1721
rect 31461 1543 31462 1721
rect 31282 0 31462 1543
use art_test  art_test_0 ~/fpga/tiny_tapeout/tt07-arond-analog/mag
timestamp 1717269366
transform 1 0 28680 0 1 5864
box -18300 -400 2000 37900
use inverter  inverter_0
timestamp 1715220266
transform 1 0 26216 0 1 2149
box 780 -1069 5116 1161
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
